module mux_mdb
  (input [15:0]  ROM_out,
   input [15:0]  RAM_out,
   input [15:0]  F_out,
   output [15:0] RAM_in,
   );

   

endmodule
