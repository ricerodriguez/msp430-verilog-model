module pipeline
  (input clk, rst);

   /*AUTOWIRE*/

   reg_file u0
     (/*AUTOINST*/);

   mux_pc u1
     (/*AUTOINST*/);
   

endmodule
