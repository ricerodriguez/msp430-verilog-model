module mux_mdb
  (// input [15:0]  MDB_out,
   // input [15:0]  CALC_out,
   // input [15:0]  F_out,
   // input [1:0]   MDB_SEL,
   // output [15:0] MDB_in,
   output [15:0] MDB_in, input [15:0] MDB_out
   );

   // Just trying to test pipeline right now
   assign MDB_in = MDB_out;
   

   

endmodule
